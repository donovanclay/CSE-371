    Mac OS X            	   2  �     �                                      ATTR      �   �  �                  �     com.apple.lastuseddate#PS         �  %com.apple.metadata:kMDItemWhereFroms   �   =  com.apple.quarantine ��%e    �    bplist00�_https://inst-fs-iad-prod.inscloudgate.net/files/19ee43c0-cac9-4551-8d74-943a75acfb96/hw3p3.sv?download=1&token=eyJ0eXAiOiJKV1QiLCJhbGciOiJIUzUxMiJ9.eyJpYXQiOjE2ODkxMzQyOTUsInVzZXJfaWQiOiIxMDAwMDAwMDQyNzM4NDIiLCJyZXNvdXJjZSI6Ii9maWxlcy8xOWVlNDNjMC1jYWM5LTQ1NTEtOGQ3NC05NDNhNzVhY2ZiOTYvaHczcDMuc3YiLCJqdGkiOiIzMzhjMzhlZi1kYjMzLTRmNzMtOTgzOC05MDQ4MDdmNWFjZTAiLCJob3N0IjoiY2FudmFzLnV3LmVkdSIsIm9yaWdpbmFsX3VybCI6Imh0dHBzOi8vYTEwLTEwNDg1OTA2NC5jbHVzdGVyMTAuY2FudmFzLXVzZXItY29udGVudC5jb20vZmlsZXMvMTA0ODU5MDY0L2Rvd25sb2FkP2Rvd25sb2FkX2ZyZD0xXHUwMDI2bm9fY2FjaGU9dHJ1ZVx1MDAyNnJlZGlyZWN0PXRydWVcdTAwMjZzZl92ZXJpZmllcj1leUowZVhBaU9pSktWMVFpTENKaGJHY2lPaUpJVXpVeE1pSjkuZXlKMWMyVnlYMmxrSWpvaU1UQXdNREF3TURBME1qY3pPRFF5SWl3aWNtOXZkRjloWTJOdmRXNTBYMmxrSWpvaU1UQXdNREF3TURBd01EZ3pPVEU1SWl3aWIyRjFkR2hmYUc5emRDSTZJbU5oYm5aaGN5NTFkeTVsWkhVaUxDSnlaWFIxY201ZmRYSnNJanB1ZFd4c0xDSm1ZV3hzWW1GamExOTFjbXdpT2lKb2RIUndjem92TDJOaGJuWmhjeTUxZHk1bFpIVXZabWxzWlhNdk1UQTBPRFU1TURZMEwyUnZkMjVzYjJGa1AyUnZkMjVzYjJGa1gyWnlaRDB4WEhVd01ESTJabUZzYkdKaFkydGZkSE05TVRZNE9URXpORE16TVNJc0ltVjRjQ0k2TVRZNE9URXpORFl6TVgwLlZaMk4wV2VYZWp0bzIyS2JBSlBMQmg5M0hVZDU1RnhKSlluczJZelBEOFFVNkFKMFpYME5FZDY5SDRpTVlUTnRfYTJPQ0xxN05yN2s4OWZpUE94V2dBIiwiZXhwIjoxNjg5MjIwNjk1fQ.fWQNOTy7bgmawOLg_NYUKFzzjWS1Xl83ynVL-YEYs7g5BIcCQP6zcQ5hZGq0u9hywQv56dABIpUY2xuSSfL5SA_?https://canvas.uw.edu/courses/1631792/files/folder/Homework/hw3  ,                           nq/0081;64ae24fc;Firefox;9494DC35-FDE9-453B-826F-7CC37ADA12D9 