    Mac OS X            	   2   �      �                                      ATTR       �   �   #                  �   #  com.apple.quarantine q/0081;650dde4c;Microsoft\x20Edge; 