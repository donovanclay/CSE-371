    Mac OS X            	   2  �     �                                      ATTR      �   �                    �   H  com.apple.macl     ,  �  %com.apple.metadata:kMDItemWhereFroms   �   =  com.apple.quarantine  ƅۗ#H����t�N��                                                      bplist00�_https://inst-fs-iad-prod.inscloudgate.net/files/e9178fff-3ef5-41be-aee9-d8af57b56640/fifo.sv?download=1&token=eyJ0eXAiOiJKV1QiLCJhbGciOiJIUzUxMiJ9.eyJpYXQiOjE2ODkxMDc5OTYsInVzZXJfaWQiOiIxMDAwMDAwMDQyNzM4NDIiLCJyZXNvdXJjZSI6Ii9maWxlcy9lOTE3OGZmZi0zZWY1LTQxYmUtYWVlOS1kOGFmNTdiNTY2NDAvZmlmby5zdiIsImp0aSI6ImE3OTIzY2Y5LTIwNWYtNDlmZC1hNzM4LTIzNDJmMjhiMWJiNiIsImhvc3QiOiJjYW52YXMudXcuZWR1Iiwib3JpZ2luYWxfdXJsIjoiaHR0cHM6Ly9hMTAtMTA0ODU5MDU4LmNsdXN0ZXIxMC5jYW52YXMtdXNlci1jb250ZW50LmNvbS9maWxlcy8xMDQ4NTkwNTgvZG93bmxvYWQ_ZG93bmxvYWRfZnJkPTFcdTAwMjZub19jYWNoZT10cnVlXHUwMDI2cmVkaXJlY3Q9dHJ1ZVx1MDAyNnNmX3ZlcmlmaWVyPWV5SjBlWEFpT2lKS1YxUWlMQ0poYkdjaU9pSklVelV4TWlKOS5leUoxYzJWeVgybGtJam9pTVRBd01EQXdNREEwTWpjek9EUXlJaXdpY205dmRGOWhZMk52ZFc1MFgybGtJam9pTVRBd01EQXdNREF3TURnek9URTVJaXdpYjJGMWRHaGZhRzl6ZENJNkltTmhiblpoY3k1MWR5NWxaSFVpTENKeVpYUjFjbTVmZFhKc0lqcHVkV3hzTENKbVlXeHNZbUZqYTE5MWNtd2lPaUpvZEhSd2N6b3ZMMk5oYm5aaGN5NTFkeTVsWkhVdlptbHNaWE12TVRBME9EVTVNRFU0TDJSdmQyNXNiMkZrUDJSdmQyNXNiMkZrWDJaeVpEMHhYSFV3TURJMlptRnNiR0poWTJ0ZmRITTlNVFk0T1RFek5ETXlPU0lzSW1WNGNDSTZNVFk0T1RFek5EWXlPWDAucl9qSEhRWkVjYThENG8xVXEzN2dBS2IwSHotMTZsdVR2VldURVhlNENxRkNpZnl3dXhJVU9odkludTdWdGg2b01mZXY0ZkJfX1poU0hfbkJxLWpnY1EiLCJleHAiOjE2ODkxOTQzOTZ9._7DA7OHJg8Sb12JayGcbdDN6L6qoqkz8IGYbbcCAFFrkVOBWR5c7wNNxDW35DlwwMNgnsVIOtORdD0yFX7FUkw_?https://canvas.uw.edu/courses/1631792/files/folder/Homework/hw3  )                           kq/0081;64ae24f9;Firefox;967C7B12-51E7-452E-A3FD-F779F925AEC6 