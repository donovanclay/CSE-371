    Mac OS X            	   2       E                                      ATTR      E    9                      com.apple.lastuseddate#PS         H  com.apple.macl     d  �  %com.apple.metadata:kMDItemWhereFroms      =  com.apple.quarantine �e    �1     ƅۗ#H����t�N��                                                      bplist00�_-https://inst-fs-iad-prod.inscloudgate.net/files/b750186e-d067-4437-8234-31334da56d36/sign_mag_add.sv?download=1&token=eyJ0eXAiOiJKV1QiLCJhbGciOiJIUzUxMiJ9.eyJpYXQiOjE2ODg1MDAwMzMsInVzZXJfaWQiOiIxMDAwMDAwMDQyNzM4NDIiLCJyZXNvdXJjZSI6Ii9maWxlcy9iNzUwMTg2ZS1kMDY3LTQ0MzctODIzNC0zMTMzNGRhNTZkMzYvc2lnbl9tYWdfYWRkLnN2IiwianRpIjoiY2YyNzgzMWEtYWYxMy00ZGQwLTg0Y2UtYjBiYTRiZjNiN2E0IiwiaG9zdCI6ImNhbnZhcy51dy5lZHUiLCJvcmlnaW5hbF91cmwiOiJodHRwczovL2ExMC0xMDQ1NjYyNTcuY2x1c3RlcjEwLmNhbnZhcy11c2VyLWNvbnRlbnQuY29tL2ZpbGVzLzEwNDU2NjI1Ny9kb3dubG9hZD9kb3dubG9hZF9mcmQ9MVx1MDAyNm5vX2NhY2hlPXRydWVcdTAwMjZyZWRpcmVjdD10cnVlXHUwMDI2c2ZfdmVyaWZpZXI9ZXlKMGVYQWlPaUpLVjFRaUxDSmhiR2NpT2lKSVV6VXhNaUo5LmV5SjFjMlZ5WDJsa0lqb2lNVEF3TURBd01EQTBNamN6T0RReUlpd2ljbTl2ZEY5aFkyTnZkVzUwWDJsa0lqb2lNVEF3TURBd01EQXdNRGd6T1RFNUlpd2liMkYxZEdoZmFHOXpkQ0k2SW1OaGJuWmhjeTUxZHk1bFpIVWlMQ0p5WlhSMWNtNWZkWEpzSWpwdWRXeHNMQ0ptWVd4c1ltRmphMTkxY213aU9pSm9kSFJ3Y3pvdkwyTmhiblpoY3k1MWR5NWxaSFV2Wm1sc1pYTXZNVEEwTlRZMk1qVTNMMlJ2ZDI1c2IyRmtQMlJ2ZDI1c2IyRmtYMlp5WkQweFhIVXdNREkyWm1Gc2JHSmhZMnRmZEhNOU1UWTRPRFV3T1RNek9TSXNJbVY0Y0NJNk1UWTRPRFV3T1RZek9YMC5FNWxiX1Bhd0szQnZGTWlDbDVfM1J1RXpyakozd2JKYjFuRDk2V3MtM3BkVHY2S05MTEV2eGx3NW9lVmZPTU5HMnZUTENTYm1kNjZPX1dIa08ydjloZyIsImV4cCI6MTY4ODU4NjQzM30.Q7HAUWEedduHKyX4nBIRCAGOYsYzzJ2xDdDEs2RRmuvA_XPBc89Nn07etkfLHR-0Dv3F-p2THCwpawvwI07P4w_?https://canvas.uw.edu/courses/1631792/files/folder/Homework/hw2  <                           ~q/0081;64a49b9c;Firefox;8334EDFB-BE11-49F4-95E5-D47DE625A490 