    Mac OS X            	   2  �                                           ATTR         �                     �   H  com.apple.macl     ,  �  %com.apple.metadata:kMDItemWhereFroms   �   =  com.apple.quarantine  ƅۗ#H����t�N��                                                      bplist00�_$https://inst-fs-iad-prod.inscloudgate.net/files/00d4a04b-ffa9-49be-b02d-a73e922d7dc5/reg_file.sv?download=1&token=eyJ0eXAiOiJKV1QiLCJhbGciOiJIUzUxMiJ9.eyJpYXQiOjE2ODkwOTk3OTMsInVzZXJfaWQiOiIxMDAwMDAwMDQyNzM4NDIiLCJyZXNvdXJjZSI6Ii9maWxlcy8wMGQ0YTA0Yi1mZmE5LTQ5YmUtYjAyZC1hNzNlOTIyZDdkYzUvcmVnX2ZpbGUuc3YiLCJqdGkiOiJmNzFjMTZlZC0xMTI1LTQwZWEtODc4Yi1lMjM1YThkNGQyNzIiLCJob3N0IjoiY2FudmFzLnV3LmVkdSIsIm9yaWdpbmFsX3VybCI6Imh0dHBzOi8vYTEwLTEwNDg1OTA2NS5jbHVzdGVyMTAuY2FudmFzLXVzZXItY29udGVudC5jb20vZmlsZXMvMTA0ODU5MDY1L2Rvd25sb2FkP2Rvd25sb2FkX2ZyZD0xXHUwMDI2bm9fY2FjaGU9dHJ1ZVx1MDAyNnJlZGlyZWN0PXRydWVcdTAwMjZzZl92ZXJpZmllcj1leUowZVhBaU9pSktWMVFpTENKaGJHY2lPaUpJVXpVeE1pSjkuZXlKMWMyVnlYMmxrSWpvaU1UQXdNREF3TURBME1qY3pPRFF5SWl3aWNtOXZkRjloWTJOdmRXNTBYMmxrSWpvaU1UQXdNREF3TURBd01EZ3pPVEU1SWl3aWIyRjFkR2hmYUc5emRDSTZJbU5oYm5aaGN5NTFkeTVsWkhVaUxDSnlaWFIxY201ZmRYSnNJanB1ZFd4c0xDSm1ZV3hzWW1GamExOTFjbXdpT2lKb2RIUndjem92TDJOaGJuWmhjeTUxZHk1bFpIVXZabWxzWlhNdk1UQTBPRFU1TURZMUwyUnZkMjVzYjJGa1AyUnZkMjVzYjJGa1gyWnlaRDB4WEhVd01ESTJabUZzYkdKaFkydGZkSE05TVRZNE9URXpORE16TkNJc0ltVjRjQ0k2TVRZNE9URXpORFl6TkgwLjd2YlJUUHYtNWk5RWctcWd1TUREM1Ezb052bDFpcjM5UkUxSVc3dUUwWS13OWYtS2FrQ3piVGw1SnBQdUtoS2VNaGFtbW13NFB3TnFEOTdEVy14S05RIiwiZXhwIjoxNjg5MTg2MTkzfQ.I-3p3kiqmZ6GRIfo-MbMvdPYaZdekOXcqvseAXBwXKU6MbDXSBPvosA4_C75DSSzM4IOekrAZTGEob_ZmmDh-Q_?https://canvas.uw.edu/courses/1631792/files/folder/Homework/hw3  3                           uq/0081;64ae24fe;Firefox;B01EF1B7-C4AA-422C-A1CE-77DF60664310 