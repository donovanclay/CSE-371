    Mac OS X            	   2       9                                      ATTR      9    -                      com.apple.lastuseddate#PS         H  com.apple.macl     d  �  %com.apple.metadata:kMDItemWhereFroms   �   =  com.apple.quarantine Q�%e    ,�+     ƅۗ#H����t�N��                                                      bplist00�_!https://inst-fs-iad-prod.inscloudgate.net/files/1638fc8c-3c85-496a-9247-d442ba42de22/fifo_tb.sv?download=1&token=eyJ0eXAiOiJKV1QiLCJhbGciOiJIUzUxMiJ9.eyJpYXQiOjE2ODkxMDk0NjMsInVzZXJfaWQiOiIxMDAwMDAwMDQyNzM4NDIiLCJyZXNvdXJjZSI6Ii9maWxlcy8xNjM4ZmM4Yy0zYzg1LTQ5NmEtOTI0Ny1kNDQyYmE0MmRlMjIvZmlmb190Yi5zdiIsImp0aSI6IjczM2UwNmZkLTRjNDQtNDNhOS05MTUzLTI4ZjJhYTdjMWQ1OSIsImhvc3QiOiJjYW52YXMudXcuZWR1Iiwib3JpZ2luYWxfdXJsIjoiaHR0cHM6Ly9hMTAtMTA0ODU5MDYzLmNsdXN0ZXIxMC5jYW52YXMtdXNlci1jb250ZW50LmNvbS9maWxlcy8xMDQ4NTkwNjMvZG93bmxvYWQ_ZG93bmxvYWRfZnJkPTFcdTAwMjZub19jYWNoZT10cnVlXHUwMDI2cmVkaXJlY3Q9dHJ1ZVx1MDAyNnNmX3ZlcmlmaWVyPWV5SjBlWEFpT2lKS1YxUWlMQ0poYkdjaU9pSklVelV4TWlKOS5leUoxYzJWeVgybGtJam9pTVRBd01EQXdNREEwTWpjek9EUXlJaXdpY205dmRGOWhZMk52ZFc1MFgybGtJam9pTVRBd01EQXdNREF3TURnek9URTVJaXdpYjJGMWRHaGZhRzl6ZENJNkltTmhiblpoY3k1MWR5NWxaSFVpTENKeVpYUjFjbTVmZFhKc0lqcHVkV3hzTENKbVlXeHNZbUZqYTE5MWNtd2lPaUpvZEhSd2N6b3ZMMk5oYm5aaGN5NTFkeTVsWkhVdlptbHNaWE12TVRBME9EVTVNRFl6TDJSdmQyNXNiMkZrUDJSdmQyNXNiMkZrWDJaeVpEMHhYSFV3TURJMlptRnNiR0poWTJ0ZmRITTlNVFk0T1RFek5ETXlOaUlzSW1WNGNDSTZNVFk0T1RFek5EWXlObjAuYktscUtwTk03VzJkYUhPSl80eDlIZVpNdXJ4dnp3RHg2XzFiS3VDdFVwX0QwcExBNTBsOXRkeXJpeEdPMzdjU0xSUGV2OWVTcmRfYjhxZlNBbTg0aVEiLCJleHAiOjE2ODkxOTU4NjN9._Ad91j047bJyIyA7_xcmrMgc-7VMdDP2txlmuwBHNDkjqnQQr79x5SZHRnCRXalKmI-yxtBH7OiJRud1yem72w_?https://canvas.uw.edu/courses/1631792/files/folder/Homework/hw3  0                           rq/0081;64ae24f7;Firefox;47DD121F-33F0-41FD-92F5-D9F3A4750137 