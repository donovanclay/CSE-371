    Mac OS X            	   2  �                                           ATTR         �  "                  �   H  com.apple.macl     ,  �  %com.apple.metadata:kMDItemWhereFroms   �   =  com.apple.quarantine  ƅۗ#H����t�N��                                                      bplist00�_&https://inst-fs-iad-prod.inscloudgate.net/files/4625c596-f4e8-4853-a112-5ac165ef567b/fifo_ctrl.sv?download=1&token=eyJ0eXAiOiJKV1QiLCJhbGciOiJIUzUxMiJ9.eyJpYXQiOjE2ODkxMzAwMzMsInVzZXJfaWQiOiIxMDAwMDAwMDQyNzM4NDIiLCJyZXNvdXJjZSI6Ii9maWxlcy80NjI1YzU5Ni1mNGU4LTQ4NTMtYTExMi01YWMxNjVlZjU2N2IvZmlmb19jdHJsLnN2IiwianRpIjoiMmY4N2RlNGEtNDMxNi00ZGZlLTljNmQtYjQ1OGQ2MGU0NDFiIiwiaG9zdCI6ImNhbnZhcy51dy5lZHUiLCJvcmlnaW5hbF91cmwiOiJodHRwczovL2ExMC0xMDQ4NTkwNjEuY2x1c3RlcjEwLmNhbnZhcy11c2VyLWNvbnRlbnQuY29tL2ZpbGVzLzEwNDg1OTA2MS9kb3dubG9hZD9kb3dubG9hZF9mcmQ9MVx1MDAyNm5vX2NhY2hlPXRydWVcdTAwMjZyZWRpcmVjdD10cnVlXHUwMDI2c2ZfdmVyaWZpZXI9ZXlKMGVYQWlPaUpLVjFRaUxDSmhiR2NpT2lKSVV6VXhNaUo5LmV5SjFjMlZ5WDJsa0lqb2lNVEF3TURBd01EQTBNamN6T0RReUlpd2ljbTl2ZEY5aFkyTnZkVzUwWDJsa0lqb2lNVEF3TURBd01EQXdNRGd6T1RFNUlpd2liMkYxZEdoZmFHOXpkQ0k2SW1OaGJuWmhjeTUxZHk1bFpIVWlMQ0p5WlhSMWNtNWZkWEpzSWpwdWRXeHNMQ0ptWVd4c1ltRmphMTkxY213aU9pSm9kSFJ3Y3pvdkwyTmhiblpoY3k1MWR5NWxaSFV2Wm1sc1pYTXZNVEEwT0RVNU1EWXhMMlJ2ZDI1c2IyRmtQMlJ2ZDI1c2IyRmtYMlp5WkQweFhIVXdNREkyWm1Gc2JHSmhZMnRmZEhNOU1UWTRPVEV6TkRNeU5DSXNJbVY0Y0NJNk1UWTRPVEV6TkRZeU5IMC4waXRzcEd6bG5vcExxZW9oQXZxbnZWcHl2a0ZXS3hpQlJpNHBoLVlnVDBmUXgwM0gzSmhIbDdfalI3Q2NPdWNVRThhZzBoNlhXZnY5Q2xLRk9GdnBDZyIsImV4cCI6MTY4OTIxNjQzM30.AL6I_4_noeTeyu1uaRwqkUrx5QqaZu29mj63to3ZGrOmY8hx9XnGpAwsedT5bxNDVbeoTAtjma8pFqQwUAfY8Q_?https://canvas.uw.edu/courses/1631792/files/folder/Homework/hw3  5                           wq/0081;64ae24f5;Firefox;114C6257-71AB-4676-B553-F0FDEDDD5343 